module slave (
    input scl,
    inout sda);
    
//------规定输入输出类型
wire scl;
wire sda;
//------规定输入输出类型

//------模块内变量定义
reg 
//------模块内变量定义

endmodule