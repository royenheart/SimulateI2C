`define idle 4'd0
`define loadDevAddr 4'd1
`define loadDevInnerAddr 4'd2
`define loadSendData 4'd3
`define sendStart 4'd4
`define sendByte 4'd5
`define recvAck 4'd6
`define verifyAck 4'd7
`define sendStop 4'd8
`define over 4'd9
