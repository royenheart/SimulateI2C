`define ridle 4'd0
`define rloadDeviceAddrFirst 4'd1
`define rloadRegisterAddr 4'd2
`define rsendStartFirst 4'd3
`define rsendByte 4'd4
`define rrecvAck 4'd5
`define rcheckAck 4'd6
`define rsendStartSecond 4'd7
`define rloadDeviceAddrSecond 4'd8
`define rreadData 4'd9
`define rrecvNotAck 4'd10
`define rclearSDA 4'd11
`define rsendStop 4'd12
`define rover 4'd13