`define idle 4'd0
`define loadDeviceAddrFirst 4'd1
`define loadRegisterAddr 4'd2
`define sendStartFirst 4'd3
`define sendByte 4'd4
`define recvAck 4'd5
`define checkAck 4'd6
`define sendStartSecond 4'd7
`define loadDeviceAddrSecond 4'd8
`define readData 4'd9
`define recvNotAck 4'd10
`define clearSDA 4'd11
`define sendStop 4'd12
`define over 4'd13